`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/19/2021 06:50:23 PM
// Design Name: 
// Module Name: graph
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module graph(
    input clk,
    input rst,
    input [100:0] init,
    output state0,
    output state1,
    output state2,
    output state3,
    output state4,
    output state5,
    output state6,
    output state7,
    output state8,
    output state9,
    output state10,
    output state11,
    output state12,
    output state13,
    output state14,
    output state15,
    output state16,
    output state17,
    output state18,
    output state19,
    output state20,
    output state21,
    output state22,
    output state23,
    output state24,
    output state25,
    output state26,
    output state27,
    output state28,
    output state29,
    output state30,
    output state31,
    output state32,
    output state33,
    output state34,
    output state35,
    output state36,
    output state37,
    output state38,
    output state39,
    output state40,
    output state41,
    output state42,
    output state43,
    output state44,
    output state45,
    output state46,
    output state47,
    output state48,
    output state49,
    output state50,
    output state51,
    output state52,
    output state53,
    output state54,
    output state55,
    output state56,
    output state57,
    output state58,
    output state59,
    output state60,
    output state61,
    output state62,
    output state63,
    output state64,
    output state65,
    output state66,
    output state67,
    output state68,
    output state69,
    output state70,
    output state71,
    output state72,
    output state73,
    output state74,
    output state75,
    output state76,
    output state77,
    output state78,
    output state79,
    output state80,
    output state81,
    output state82,
    output state83,
    output state84,
    output state85,
    output state86,
    output state87,
    output state88,
    output state89,
    output state90,
    output state91,
    output state92,
    output state93,
    output state94,
    output state95,
    output state96,
    output state97,
    output state98,
    output state99
    );


    reg out0;
    reg out1; 
    reg out3;
    reg out4;
    reg out5;
    reg out6;
    reg out7;
    reg out8;
    reg out9;
    reg out10;
    reg out11;
    reg out12;
    reg out13;
    reg out14;
    reg out15;
    reg out16;
    reg out17;
    reg out18;
    reg out19;
    reg out20;
    reg out21;
    reg out22;
    reg out23;
    reg out24;
    reg out25;
    reg out26;
    reg out27;
    reg out28;
    reg out29;
    reg out30;
    reg out31;
    reg out32;
    reg out33;
    reg out34;
    reg out35;
    reg out36;
    reg out37;
    reg out38;
    reg out39;
    reg out40;
    reg out41;
    reg out42;
    reg out43;
    reg out44;
    reg out45;
    reg out46;
    reg out47;
    reg out48;
    reg out49;
    reg out50;
    reg out51;
    reg out52;
    reg out53;
    reg out54;
    reg out55;
    reg out56;
    reg out57;
    reg out58;
    reg out59;
    reg out60;
    reg out61;
    reg out62;
    reg out63;
    reg out64;
    reg out65;
    reg out66;
    reg out67;
    reg out68;
    reg out69;
    reg out70;
    reg out71;
    reg out72;
    reg out73;
    reg out74;
    reg out75;
    reg out76;
    reg out77;
    reg out78;
    reg out79;
    reg out80;
    reg out81;
    reg out82;
    reg out83;
    reg out84;
    reg out85;
    reg out86;
    reg out87;
    reg out88;
    reg out89;
    reg out90;
    reg out91;
    reg out92;
    reg out93;
    reg out94;
    reg out95;
    reg out96;
    reg out97;
    reg out98;
    reg out99;
    reg out100;
    reg out101;
    reg out102;
    reg out103;
    reg out104;
    reg out105;
    reg out106;
    reg out107;
    reg out108;
    reg out109;
    reg out110;
    reg out111;
    reg out112;
    reg out113;
    reg out114;
    reg out115;
    reg out116;
    reg out117;
    reg out118;
    reg out119;
    reg out120;
    reg out121;
    reg out122;
    reg out123;
    reg out124;
    reg out125;
    reg out126;
    reg out127;
    reg out128;
    reg out129;
    reg out130;
    reg out131;
    reg out132;
    reg out133;
    reg out134;
    reg out135;
    reg out136;
    reg out137;
    reg out138;
    reg out139;
    reg out140;
    reg out141;
    reg out142;
    reg out143;

    CELL cell_0(clk, rst, init[0], 1'b0, out1, out12, 1'b0, out0);
    CELL cell_1(clk, rst, init[1], 1'b0, out2, out13, out0, out1);
    CELL cell_2(clk, rst, init[2], 1'b0, out3, out14, out1, out2);
    CELL cell_3(clk, rst, init[3], 1'b0, out4, out15, out2, out3);
    CELL cell_4(clk, rst, init[4], 1'b0, out5, out16, out3, out4);
    CELL cell_5(clk, rst, init[5], 1'b0, out6, out17, out4, out5);
    CELL cell_6(clk, rst, init[6], 1'b0, out7, out18, out5, out6);
    CELL cell_7(clk, rst, init[7], 1'b0, out8, out19, out6, out7);
    CELL cell_8(clk, rst, init[8], 1'b0, out9, out20, out7, out8);
    CELL cell_9(clk, rst, init[9], 1'b0, out10, out21, out8, out9);
    CELL cell_10(clk, rst, init[10], 1'b0, out11, out22, out9, out10);
    CELL cell_11(clk, rst, init[11], 1'b0, 1'b0, out23, out10, out11);
    CELL cell_12(clk, rst, init[12], out0, out13, out24, 1'b0, out12);
    CELL cell_13(clk, rst, init[13], out1, out14, out25, out12, out13);
    CELL cell_14(clk, rst, init[14], out2, out15, out26, out13, out14);
    CELL cell_15(clk, rst, init[15], out3, out16, out27, out14, out15);
    CELL cell_16(clk, rst, init[16], out4, out17, out28, out15, out16);
    CELL cell_17(clk, rst, init[17], out5, out18, out29, out16, out17);
    CELL cell_18(clk, rst, init[18], out6, out19, out30, out17, out18);
    CELL cell_19(clk, rst, init[19], out7, out20, out31, out18, out19);
    CELL cell_20(clk, rst, init[20], out8, out21, out32, out19, out20);
    CELL cell_21(clk, rst, init[21], out9, out22, out33, out20, out21);
    CELL cell_22(clk, rst, init[22], out10, out23, out34, out21, out22);
    CELL cell_23(clk, rst, init[23], out11, 1'b0, out35, out22, out23);
    CELL cell_24(clk, rst, init[24], out12, out25, out36, 1'b0, out24);
    CELL cell_25(clk, rst, init[25], out13, out26, out37, out24, out25);
    CELL cell_26(clk, rst, init[26], out14, out27, out38, out25, out26);
    CELL cell_27(clk, rst, init[27], out15, out28, out39, out26, out27);
    CELL cell_28(clk, rst, init[28], out16, out29, out40, out27, out28);
    CELL cell_29(clk, rst, init[29], out17, out30, out41, out28, out29);
    CELL cell_30(clk, rst, init[30], out18, out31, out42, out29, out30);
    CELL cell_31(clk, rst, init[31], out19, out32, out43, out30, out31);
    CELL cell_32(clk, rst, init[32], out20, out33, out44, out31, out32);
    CELL cell_33(clk, rst, init[33], out21, out34, out45, out32, out33);
    CELL cell_34(clk, rst, init[34], out22, out35, out46, out33, out34);
    CELL cell_35(clk, rst, init[35], out23, 1'b0, out47, out34, out35);
    CELL cell_36(clk, rst, init[36], out24, out37, out48, 1'b0, out36);
    CELL cell_37(clk, rst, init[37], out25, out38, out49, out36, out37);
    CELL cell_38(clk, rst, init[38], out26, out39, out50, out37, out38);
    CELL cell_39(clk, rst, init[39], out27, out40, out51, out38, out39);
    CELL cell_40(clk, rst, init[40], out28, out41, out52, out39, out40);
    CELL cell_41(clk, rst, init[41], out29, out42, out53, out40, out41);
    CELL cell_42(clk, rst, init[42], out30, out43, out54, out41, out42);
    CELL cell_43(clk, rst, init[43], out31, out44, out55, out42, out43);
    CELL cell_44(clk, rst, init[44], out32, out45, out56, out43, out44);
    CELL cell_45(clk, rst, init[45], out33, out46, out57, out44, out45);
    CELL cell_46(clk, rst, init[46], out34, out47, out58, out45, out46);
    CELL cell_47(clk, rst, init[47], out35, 1'b0, out59, out46, out47);
    CELL cell_48(clk, rst, init[48], out36, out49, out60, 1'b0, out48);
    CELL cell_49(clk, rst, init[49], out37, out50, out61, out48, out49);
    CELL cell_50(clk, rst, init[50], out38, out51, out62, out49, out50);
    CELL cell_51(clk, rst, init[51], out39, out52, out63, out50, out51);
    CELL cell_52(clk, rst, init[52], out40, out53, out64, out51, out52);
    CELL cell_53(clk, rst, init[53], out41, out54, out65, out52, out53);
    CELL cell_54(clk, rst, init[54], out42, out55, out66, out53, out54);
    CELL cell_55(clk, rst, init[55], out43, out56, out67, out54, out55);
    CELL cell_56(clk, rst, init[56], out44, out57, out68, out55, out56);
    CELL cell_57(clk, rst, init[57], out45, out58, out69, out56, out57);
    CELL cell_58(clk, rst, init[58], out46, out59, out70, out57, out58);
    CELL cell_59(clk, rst, init[59], out47, 1'b0, out71, out58, out59);
    CELL cell_60(clk, rst, init[60], out48, out61, out72, 1'b0, out60);
    CELL cell_61(clk, rst, init[61], out49, out62, out73, out60, out61);
    CELL cell_62(clk, rst, init[62], out50, out63, out74, out61, out62);
    CELL cell_63(clk, rst, init[63], out51, out64, out75, out62, out63);
    CELL cell_64(clk, rst, init[64], out52, out65, out76, out63, out64);
    CELL cell_65(clk, rst, init[65], out53, out66, out77, out64, out65);
    CELL cell_66(clk, rst, init[66], out54, out67, out78, out65, out66);
    CELL cell_67(clk, rst, init[67], out55, out68, out79, out66, out67);
    CELL cell_68(clk, rst, init[68], out56, out69, out80, out67, out68);
    CELL cell_69(clk, rst, init[69], out57, out70, out81, out68, out69);
    CELL cell_70(clk, rst, init[70], out58, out71, out82, out69, out70);
    CELL cell_71(clk, rst, init[71], out59, 1'b0, out83, out70, out71);
    CELL cell_72(clk, rst, init[72], out60, out73, out84, 1'b0, out72);
    CELL cell_73(clk, rst, init[73], out61, out74, out85, out72, out73);
    CELL cell_74(clk, rst, init[74], out62, out75, out86, out73, out74);
    CELL cell_75(clk, rst, init[75], out63, out76, out87, out74, out75);
    CELL cell_76(clk, rst, init[76], out64, out77, out88, out75, out76);
    CELL cell_77(clk, rst, init[77], out65, out78, out89, out76, out77);
    CELL cell_78(clk, rst, init[78], out66, out79, out90, out77, out78);
    CELL cell_79(clk, rst, init[79], out67, out80, out91, out78, out79);
    CELL cell_80(clk, rst, init[80], out68, out81, out92, out79, out80);
    CELL cell_81(clk, rst, init[81], out69, out82, out93, out80, out81);
    CELL cell_82(clk, rst, init[82], out70, out83, out94, out81, out82);
    CELL cell_83(clk, rst, init[83], out71, 1'b0, out95, out82, out83);
    CELL cell_84(clk, rst, init[84], out72, out85, out96, 1'b0, out84);
    CELL cell_85(clk, rst, init[85], out73, out86, out97, out84, out85);
    CELL cell_86(clk, rst, init[86], out74, out87, out98, out85, out86);
    CELL cell_87(clk, rst, init[87], out75, out88, out99, out86, out87);
    CELL cell_88(clk, rst, init[88], out76, out89, out100, out87, out88);
    CELL cell_89(clk, rst, init[89], out77, out90, out101, out88, out89);
    CELL cell_90(clk, rst, init[90], out78, out91, out102, out89, out90);
    CELL cell_91(clk, rst, init[91], out79, out92, out103, out90, out91);
    CELL cell_92(clk, rst, init[92], out80, out93, out104, out91, out92);
    CELL cell_93(clk, rst, init[93], out81, out94, out105, out92, out93);
    CELL cell_94(clk, rst, init[94], out82, out95, out106, out93, out94);
    CELL cell_95(clk, rst, init[95], out83, 1'b0, out107, out94, out95);
    CELL cell_96(clk, rst, init[96], out84, out97, out108, 1'b0, out96);
    CELL cell_97(clk, rst, init[97], out85, out98, out109, out96, out97);
    CELL cell_98(clk, rst, init[98], out86, out99, out110, out97, out98);
    CELL cell_99(clk, rst, init[99], out87, out100, out111, out98, out99);
    CELL cell_100(clk, rst, init[100], out88, out101, out112, out99, out100);
    CELL cell_101(clk, rst, init[101], out89, out102, out113, out100, out101);
    CELL cell_102(clk, rst, init[102], out90, out103, out114, out101, out102);
    CELL cell_103(clk, rst, init[103], out91, out104, out115, out102, out103);
    CELL cell_104(clk, rst, init[104], out92, out105, out116, out103, out104);
    CELL cell_105(clk, rst, init[105], out93, out106, out117, out104, out105);
    CELL cell_106(clk, rst, init[106], out94, out107, out118, out105, out106);
    CELL cell_107(clk, rst, init[107], out95, 1'b0, out119, out106, out107);
    CELL cell_108(clk, rst, init[108], out96, out109, out120, 1'b0, out108);
    CELL cell_109(clk, rst, init[109], out97, out110, out121, out108, out109);
    CELL cell_110(clk, rst, init[110], out98, out111, out122, out109, out110);
    CELL cell_111(clk, rst, init[111], out99, out112, out123, out110, out111);
    CELL cell_112(clk, rst, init[112], out100, out113, out124, out111, out112);
    CELL cell_113(clk, rst, init[113], out101, out114, out125, out112, out113);
    CELL cell_114(clk, rst, init[114], out102, out115, out126, out113, out114);
    CELL cell_115(clk, rst, init[115], out103, out116, out127, out114, out115);
    CELL cell_116(clk, rst, init[116], out104, out117, out128, out115, out116);
    CELL cell_117(clk, rst, init[117], out105, out118, out129, out116, out117);
    CELL cell_118(clk, rst, init[118], out106, out119, out130, out117, out118);
    CELL cell_119(clk, rst, init[119], out107, 1'b0, out131, out118, out119);
    CELL cell_120(clk, rst, init[120], out108, out121, out132, 1'b0, out120);
    CELL cell_121(clk, rst, init[121], out109, out122, out133, out120, out121);
    CELL cell_122(clk, rst, init[122], out110, out123, out134, out121, out122);
    CELL cell_123(clk, rst, init[123], out111, out124, out135, out122, out123);
    CELL cell_124(clk, rst, init[124], out112, out125, out136, out123, out124);
    CELL cell_125(clk, rst, init[125], out113, out126, out137, out124, out125);
    CELL cell_126(clk, rst, init[126], out114, out127, out138, out125, out126);
    CELL cell_127(clk, rst, init[127], out115, out128, out139, out126, out127);
    CELL cell_128(clk, rst, init[128], out116, out129, out140, out127, out128);
    CELL cell_129(clk, rst, init[129], out117, out130, out141, out128, out129);
    CELL cell_130(clk, rst, init[130], out118, out131, out142, out129, out130);
    CELL cell_131(clk, rst, init[131], out119, 1'b0, out143, out130, out131);
    CELL cell_132(clk, rst, init[132], out120, out133, 1'b0, 1'b0, out132);
    CELL cell_133(clk, rst, init[133], out121, out134, 1'b0, out132, out133);
    CELL cell_134(clk, rst, init[134], out122, out135, 1'b0, out133, out134);
    CELL cell_135(clk, rst, init[135], out123, out136, 1'b0, out134, out135);
    CELL cell_136(clk, rst, init[136], out124, out137, 1'b0, out135, out136);
    CELL cell_137(clk, rst, init[137], out125, out138, 1'b0, out136, out137);
    CELL cell_138(clk, rst, init[138], out126, out139, 1'b0, out137, out138);
    CELL cell_139(clk, rst, init[139], out127, out140, 1'b0, out138, out139);
    CELL cell_140(clk, rst, init[140], out128, out141, 1'b0, out139, out140);
    CELL cell_141(clk, rst, init[141], out129, out142, 1'b0, out140, out141);
    CELL cell_142(clk, rst, init[142], out130, out143, 1'b0, out141, out142);
    CELL cell_143(clk, rst, init[143], out131, 1'b0, 1'b0, out142, out143);

    assign state0 = out13;
    assign state1 = out14;
    assign state2 = out15;
    assign state3 = out16;
    assign state4 = out17;
    assign state5 = out18;
    assign state6 = out19;
    assign state7 = out20;
    assign state8 = out21;
    assign state9 = out22;
    assign state10 = out25;
    assign state11 = out26;
    assign state12 = out27;
    assign state13 = out28;
    assign state14 = out29;
    assign state15 = out30;
    assign state16 = out31;
    assign state17 = out32;
    assign state18 = out33;
    assign state19 = out34;
    assign state20 = out37;
    assign state21 = out38;
    assign state22 = out39;
    assign state23 = out40;
    assign state24 = out41;
    assign state25 = out42;
    assign state26 = out43;
    assign state27 = out44;
    assign state28 = out45;
    assign state29 = out46;
    assign state30 = out49;
    assign state31 = out50;
    assign state32 = out51;
    assign state33 = out52;
    assign state34 = out53;
    assign state35 = out54;
    assign state36 = out55;
    assign state37 = out56;
    assign state38 = out57;
    assign state39 = out58;
    assign state40 = out61;
    assign state41 = out62;
    assign state42 = out63;
    assign state43 = out64;
    assign state44 = out65;
    assign state45 = out66;
    assign state46 = out67;
    assign state47 = out68;
    assign state48 = out69;
    assign state49 = out70;
    assign state50 = out73;
    assign state51 = out74;
    assign state52 = out75;
    assign state53 = out76;
    assign state54 = out77;
    assign state55 = out78;
    assign state56 = out79;
    assign state57 = out80;
    assign state58 = out81;
    assign state59 = out82;
    assign state60 = out85;
    assign state61 = out86;
    assign state62 = out87;
    assign state63 = out88;
    assign state64 = out89;
    assign state65 = out90;
    assign state66 = out91;
    assign state67 = out92;
    assign state68 = out93;
    assign state69 = out94;
    assign state70 = out97;
    assign state71 = out98;
    assign state72 = out99;
    assign state73 = out100;
    assign state74 = out101;
    assign state75 = out102;
    assign state76 = out103;
    assign state77 = out104;
    assign state78 = out105;
    assign state79 = out106;
    assign state80 = out109;
    assign state81 = out110;
    assign state82 = out111;
    assign state83 = out112;
    assign state84 = out113;
    assign state85 = out114;
    assign state86 = out115;
    assign state87 = out116;
    assign state88 = out117;
    assign state89 = out118;
    assign state90 = out121;
    assign state91 = out122;
    assign state92 = out123;
    assign state93 = out124;
    assign state94 = out125;
    assign state95 = out126;
    assign state96 = out127;
    assign state97 = out128;
    assign state98 = out129;
    assign state99 = out130;

endmodule